LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

USE work.aes_pkg.ALL;

ENTITY sbox IS
    PORT (
        input_byte  : IN  byte_t;
        output_byte : OUT byte_t
    );
END sbox;

ARCHITECTURE Behaviour OF sbox IS
BEGIN
    WITH input_byte SELECT output_byte <=
        -- Row 0x00 - 0x0F                                                                                                                                                                  
        x"63" WHEN x"00", x"7C" WHEN x"01", x"77" WHEN x"02", x"7B" WHEN x"03",
        x"F2" WHEN x"04", x"6B" WHEN x"05", x"6F" WHEN x"06", x"C5" WHEN x"07",
        x"30" WHEN x"08", x"01" WHEN x"09", x"67" WHEN x"0A", x"2B" WHEN x"0B",
        x"FE" WHEN x"0C", x"D7" WHEN x"0D", x"AB" WHEN x"0E", x"76" WHEN x"0F",
        -- Row 0x10 - 0x1F                                                                                                                                                                  
        x"CA" WHEN x"10", x"82" WHEN x"11", x"C9" WHEN x"12", x"7D" WHEN x"13",
        x"FA" WHEN x"14", x"59" WHEN x"15", x"47" WHEN x"16", x"F0" WHEN x"17",
        x"AD" WHEN x"18", x"D4" WHEN x"19", x"A2" WHEN x"1A", x"AF" WHEN x"1B",
        x"9C" WHEN x"1C", x"A4" WHEN x"1D", x"72" WHEN x"1E", x"C0" WHEN x"1F",
        -- Row 0x20 - 0x2F                                                                                                                                                                  
        x"B7" WHEN x"20", x"FD" WHEN x"21", x"93" WHEN x"22", x"26" WHEN x"23",
        x"36" WHEN x"24", x"3F" WHEN x"25", x"F7" WHEN x"26", x"CC" WHEN x"27",
        x"34" WHEN x"28", x"A5" WHEN x"29", x"E5" WHEN x"2A", x"F1" WHEN x"2B",
        x"71" WHEN x"2C", x"D8" WHEN x"2D", x"31" WHEN x"2E", x"15" WHEN x"2F",
        -- Row 0x30 - 0x3F                                                                                                                                                                  
        x"04" WHEN x"30", x"C7" WHEN x"31", x"23" WHEN x"32", x"C3" WHEN x"33",
        x"18" WHEN x"34", x"96" WHEN x"35", x"05" WHEN x"36", x"9A" WHEN x"37",
        x"07" WHEN x"38", x"12" WHEN x"39", x"80" WHEN x"3A", x"E2" WHEN x"3B",
        x"EB" WHEN x"3C", x"27" WHEN x"3D", x"B2" WHEN x"3E", x"75" WHEN x"3F",
        -- Row 0x40 - 0x4F                                                                                                                                                                  
        x"09" WHEN x"40", x"83" WHEN x"41", x"2C" WHEN x"42", x"1A" WHEN x"43",
        x"1B" WHEN x"44", x"6E" WHEN x"45", x"5A" WHEN x"46", x"A0" WHEN x"47",
        x"52" WHEN x"48", x"3B" WHEN x"49", x"D6" WHEN x"4A", x"B3" WHEN x"4B",
        x"29" WHEN x"4C", x"E3" WHEN x"4D", x"2F" WHEN x"4E", x"84" WHEN x"4F",
        -- Row 0x50 - 0x5F                                                                                                                                                                  
        x"53" WHEN x"50", x"D1" WHEN x"51", x"00" WHEN x"52", x"ED" WHEN x"53",
        x"20" WHEN x"54", x"FC" WHEN x"55", x"B1" WHEN x"56", x"5B" WHEN x"57",
        x"6A" WHEN x"58", x"CB" WHEN x"59", x"BE" WHEN x"5A", x"39" WHEN x"5B",
        x"4A" WHEN x"5C", x"4C" WHEN x"5D", x"58" WHEN x"5E", x"CF" WHEN x"5F",
        -- Row 0x60 - 0x6F                                                                                                                                                                  
        x"D0" WHEN x"60", x"EF" WHEN x"61", x"AA" WHEN x"62", x"FB" WHEN x"63",
        x"43" WHEN x"64", x"4D" WHEN x"65", x"33" WHEN x"66", x"85" WHEN x"67",
        x"45" WHEN x"68", x"F9" WHEN x"69", x"02" WHEN x"6A", x"7F" WHEN x"6B",
        x"50" WHEN x"6C", x"3C" WHEN x"6D", x"9F" WHEN x"6E", x"A8" WHEN x"6F",
        -- Row 0x70 - 0x7F                                                                                                                                                                  
        x"51" WHEN x"70", x"A3" WHEN x"71", x"40" WHEN x"72", x"8F" WHEN x"73",
        x"92" WHEN x"74", x"9D" WHEN x"75", x"38" WHEN x"76", x"F5" WHEN x"77",
        x"BC" WHEN x"78", x"B6" WHEN x"79", x"DA" WHEN x"7A", x"21" WHEN x"7B",
        x"10" WHEN x"7C", x"FF" WHEN x"7D", x"F3" WHEN x"7E", x"D2" WHEN x"7F",
        -- Row 0x80 - 0x8F                                                                                                                                                                  
        x"CD" WHEN x"80", x"0C" WHEN x"81", x"13" WHEN x"82", x"EC" WHEN x"83",
        x"5F" WHEN x"84", x"97" WHEN x"85", x"44" WHEN x"86", x"17" WHEN x"87",
        x"C4" WHEN x"88", x"A7" WHEN x"89", x"7E" WHEN x"8A", x"3D" WHEN x"8B",
        x"64" WHEN x"8C", x"5D" WHEN x"8D", x"19" WHEN x"8E", x"73" WHEN x"8F",
        -- Row 0x90 - 0x9F                                                                                                                                                                  
        x"60" WHEN x"90", x"81" WHEN x"91", x"4F" WHEN x"92", x"DC" WHEN x"93",
        x"22" WHEN x"94", x"2A" WHEN x"95", x"90" WHEN x"96", x"88" WHEN x"97",
        x"46" WHEN x"98", x"EE" WHEN x"99", x"B8" WHEN x"9A", x"14" WHEN x"9B",
        x"DE" WHEN x"9C", x"5E" WHEN x"9D", x"0B" WHEN x"9E", x"DB" WHEN x"9F",
        -- Row 0xA0 - 0xAF                                                                                                                                                                  
        x"E0" WHEN x"A0", x"32" WHEN x"A1", x"3A" WHEN x"A2", x"0A" WHEN x"A3",
        x"49" WHEN x"A4", x"06" WHEN x"A5", x"24" WHEN x"A6", x"5C" WHEN x"A7",
        x"C2" WHEN x"A8", x"D3" WHEN x"A9", x"AC" WHEN x"AA", x"62" WHEN x"AB",
        x"91" WHEN x"AC", x"95" WHEN x"AD", x"E4" WHEN x"AE", x"79" WHEN x"AF",
        -- Row 0xB0 - 0xBF                                                                                                                                                                  
        x"E7" WHEN x"B0", x"C8" WHEN x"B1", x"37" WHEN x"B2", x"6D" WHEN x"B3",
        x"8D" WHEN x"B4", x"D5" WHEN x"B5", x"4E" WHEN x"B6", x"A9" WHEN x"B7",
        x"6C" WHEN x"B8", x"56" WHEN x"B9", x"F4" WHEN x"BA", x"EA" WHEN x"BB",
        x"65" WHEN x"BC", x"7A" WHEN x"BD", x"AE" WHEN x"BE", x"08" WHEN x"BF",
        -- Row 0xC0 - 0xCF                                                                                                                                                                  
        x"BA" WHEN x"C0", x"78" WHEN x"C1", x"25" WHEN x"C2", x"2E" WHEN x"C3",
        x"1C" WHEN x"C4", x"A6" WHEN x"C5", x"B4" WHEN x"C6", x"C6" WHEN x"C7",
        x"E8" WHEN x"C8", x"DD" WHEN x"C9", x"74" WHEN x"CA", x"1F" WHEN x"CB",
        x"4B" WHEN x"CC", x"BD" WHEN x"CD", x"8B" WHEN x"CE", x"8A" WHEN x"CF",
        -- Row 0xD0 - 0xDF                                                                                                                                                                  
        x"70" WHEN x"D0", x"3E" WHEN x"D1", x"B5" WHEN x"D2", x"66" WHEN x"D3",
        x"48" WHEN x"D4", x"03" WHEN x"D5", x"F6" WHEN x"D6", x"0E" WHEN x"D7",
        x"61" WHEN x"D8", x"35" WHEN x"D9", x"57" WHEN x"DA", x"B9" WHEN x"DB",
        x"86" WHEN x"DC", x"C1" WHEN x"DD", x"1D" WHEN x"DE", x"9E" WHEN x"DF",
        -- Row 0xE0 - 0xEF                                                                                                                                                                  
        x"E1" WHEN x"E0", x"F8" WHEN x"E1", x"98" WHEN x"E2", x"11" WHEN x"E3",
        x"69" WHEN x"E4", x"D9" WHEN x"E5", x"8E" WHEN x"E6", x"94" WHEN x"E7",
        x"9B" WHEN x"E8", x"1E" WHEN x"E9", x"87" WHEN x"EA", x"E9" WHEN x"EB",
        x"CE" WHEN x"EC", x"55" WHEN x"ED", x"28" WHEN x"EE", x"DF" WHEN x"EF",
        -- Row 0xF0 - 0xFF                                                                                                                                                                  
        x"8C" WHEN x"F0", x"A1" WHEN x"F1", x"89" WHEN x"F2", x"0D" WHEN x"F3",
        x"BF" WHEN x"F4", x"E6" WHEN x"F5", x"42" WHEN x"F6", x"68" WHEN x"F7",
        x"41" WHEN x"F8", x"99" WHEN x"F9", x"2D" WHEN x"FA", x"0F" WHEN x"FB",
        x"B0" WHEN x"FC", x"54" WHEN x"FD", x"BB" WHEN x"FE", x"16" WHEN x"FF",
        -- should never happen :)                                                                                                                                                    
        x"00" WHEN OTHERS;
END Behaviour;